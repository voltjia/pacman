	component pacman_soc is
		port (
			clk_clk          : in    std_logic                     := 'X';             -- clk
			gpio_0_in_port   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- in_port
			gpio_0_out_port  : out   std_logic_vector(31 downto 0);                    -- out_port
			gpio_1_in_port   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- in_port
			gpio_1_out_port  : out   std_logic_vector(31 downto 0);                    -- out_port
			gpio_2_in_port   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- in_port
			gpio_2_out_port  : out   std_logic_vector(31 downto 0);                    -- out_port
			gpio_3_in_port   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- in_port
			gpio_3_out_port  : out   std_logic_vector(31 downto 0);                    -- out_port
			reset_reset_n    : in    std_logic                     := 'X';             -- reset_n
			sdram_clk_clk    : out   std_logic;                                        -- clk
			sdram_wire_addr  : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_wire_ba    : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_wire_cas_n : out   std_logic;                                        -- cas_n
			sdram_wire_cke   : out   std_logic;                                        -- cke
			sdram_wire_cs_n  : out   std_logic;                                        -- cs_n
			sdram_wire_dq    : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_wire_dqm   : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_wire_ras_n : out   std_logic;                                        -- ras_n
			sdram_wire_we_n  : out   std_logic;                                        -- we_n
			spi_MISO         : in    std_logic                     := 'X';             -- MISO
			spi_MOSI         : out   std_logic;                                        -- MOSI
			spi_SCLK         : out   std_logic;                                        -- SCLK
			spi_SS_n         : out   std_logic;                                        -- SS_n
			usb_gpx_export   : in    std_logic                     := 'X';             -- export
			usb_irq_export   : in    std_logic                     := 'X';             -- export
			usb_rst_export   : out   std_logic;                                        -- export
			control_export   : out   std_logic_vector(31 downto 0)                     -- export
		);
	end component pacman_soc;

	u0 : component pacman_soc
		port map (
			clk_clk          => CONNECTED_TO_clk_clk,          --        clk.clk
			gpio_0_in_port   => CONNECTED_TO_gpio_0_in_port,   --     gpio_0.in_port
			gpio_0_out_port  => CONNECTED_TO_gpio_0_out_port,  --           .out_port
			gpio_1_in_port   => CONNECTED_TO_gpio_1_in_port,   --     gpio_1.in_port
			gpio_1_out_port  => CONNECTED_TO_gpio_1_out_port,  --           .out_port
			gpio_2_in_port   => CONNECTED_TO_gpio_2_in_port,   --     gpio_2.in_port
			gpio_2_out_port  => CONNECTED_TO_gpio_2_out_port,  --           .out_port
			gpio_3_in_port   => CONNECTED_TO_gpio_3_in_port,   --     gpio_3.in_port
			gpio_3_out_port  => CONNECTED_TO_gpio_3_out_port,  --           .out_port
			reset_reset_n    => CONNECTED_TO_reset_reset_n,    --      reset.reset_n
			sdram_clk_clk    => CONNECTED_TO_sdram_clk_clk,    --  sdram_clk.clk
			sdram_wire_addr  => CONNECTED_TO_sdram_wire_addr,  -- sdram_wire.addr
			sdram_wire_ba    => CONNECTED_TO_sdram_wire_ba,    --           .ba
			sdram_wire_cas_n => CONNECTED_TO_sdram_wire_cas_n, --           .cas_n
			sdram_wire_cke   => CONNECTED_TO_sdram_wire_cke,   --           .cke
			sdram_wire_cs_n  => CONNECTED_TO_sdram_wire_cs_n,  --           .cs_n
			sdram_wire_dq    => CONNECTED_TO_sdram_wire_dq,    --           .dq
			sdram_wire_dqm   => CONNECTED_TO_sdram_wire_dqm,   --           .dqm
			sdram_wire_ras_n => CONNECTED_TO_sdram_wire_ras_n, --           .ras_n
			sdram_wire_we_n  => CONNECTED_TO_sdram_wire_we_n,  --           .we_n
			spi_MISO         => CONNECTED_TO_spi_MISO,         --        spi.MISO
			spi_MOSI         => CONNECTED_TO_spi_MOSI,         --           .MOSI
			spi_SCLK         => CONNECTED_TO_spi_SCLK,         --           .SCLK
			spi_SS_n         => CONNECTED_TO_spi_SS_n,         --           .SS_n
			usb_gpx_export   => CONNECTED_TO_usb_gpx_export,   --    usb_gpx.export
			usb_irq_export   => CONNECTED_TO_usb_irq_export,   --    usb_irq.export
			usb_rst_export   => CONNECTED_TO_usb_rst_export,   --    usb_rst.export
			control_export   => CONNECTED_TO_control_export    --    control.export
		);

